library ieee;
use ieee.std_logic_1164.all;
---------------------------------
entity vote5 is
    port
    (   a  : in  std_logic_vector(4 downto 0);
        f  : out std_logic );
end;
---------------------------------
architecture arch of vote5 is
begin
    -- add your code below
end architecture;

