LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- ʵ�嶨�壺song
-- ���ڸ��ݵ�ǰ������� (music_num) �����Ӧ�������ź� (tone2)
ENTITY song IS
	PORT (
		clk8hz : IN STD_LOGIC; -- ���� 8Hz ʱ���ź�
		tone2 : OUT INTEGER RANGE 0 TO 10; -- ��������ź�
		music_num : IN INTEGER RANGE 0 TO 2 := 0 -- ��ǰ������� (Ĭ��Ϊ 0)
	);
END ENTITY;

ARCHITECTURE song_arch OF song IS
	-- �ڲ��źŶ���
	SIGNAL ptr1 : INTEGER RANGE 0 TO 239; -- little_star ��Ŀָ��
	SIGNAL ptr2 : INTEGER RANGE 0 TO 181; -- thx ��Ŀָ��
	SIGNAL ptr3 : INTEGER RANGE 0 TO 264;
	SIGNAL mn_former : INTEGER RANGE 0 TO 2 := 0; -- ��¼��һ�������, �����и���

	-- ����������������������
	TYPE pitch_array1 IS ARRAY (0 TO 239) OF INTEGER; -- ��Ŀ 1 ����������
	TYPE pitch_array2 IS ARRAY (0 TO 181) OF INTEGER; -- ��Ŀ 2 ����������
	TYPE pitch_array3 IS ARRAY (0 TO 255) OF INTEGER; -- ��Ŀ 3 ����������

	-- ��Ŀ 1��С���ǵ���������
	CONSTANT little_star : pitch_array1 := (
		1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 5, 5, 5, 5, 0, 5, 5, 5, 5, 0, 6, 6, 6, 6, 0, 6, 6, 6, 6, 0,
		5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 3, 3, 3, 3, 0, 3, 3, 3, 3, 0,
		2, 2, 2, 2, 0, 2, 2, 2, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 5, 5, 5, 5, 0, 5, 5, 5, 5, 0,
		4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 3, 3, 3, 3, 0, 3, 3, 3, 3, 0, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0,
		5, 5, 5, 5, 0, 5, 5, 5, 5, 0, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 3, 3, 3, 3, 0, 3, 3, 3, 3, 0,
		2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 5, 5, 5, 5, 0, 5, 5, 5, 5, 0,
		6, 6, 6, 6, 0, 6, 6, 6, 6, 0, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0,
		3, 3, 3, 3, 0, 3, 3, 3, 3, 0, 2, 2, 2, 2, 0, 2, 2, 2, 2, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0
	);

	-- ��Ŀ 2����л����������������
	CONSTANT thx : pitch_array2 := (
		4, 4, 0, 5, 5, 0, 6, 6, 0, 8, 8, 0, 6, 6, 0, 6, 6, 6, 6, 0, 5, 0, 5, 4, 4, 0, 5, 5, 5, 5,
		0, 4, 4, 0, 2, 2, 0, 4, 4, 0, 5, 5, 0, 6, 6, 6, 6, 6, 6, 6, 6, 0, 4, 4, 0, 2, 2, 0, 4, 4,
		4, 4, 0, 1, 0, 1, 5, 5, 0, 4, 4, 4, 4, 0, 6, 6, 0, 5, 5, 0, 5, 5, 0, 4, 4, 0, 5, 5, 5, 5,
		0, 4, 4, 0, 5, 5, 0, 6, 6, 0, 8, 8, 0, 6, 6, 0, 6, 6, 6, 6, 0, 5, 0, 5, 4, 4, 0, 5, 5, 5,
		5, 0, 4, 4, 0, 2, 2, 0, 4, 4, 0, 5, 5, 0, 6, 6, 6, 6, 6, 6, 6, 6, 0, 4, 4, 0, 2, 2, 0, 4,
		4, 4, 4, 0, 1, 0, 1, 5, 5, 0, 4, 4, 4, 4, 0, 6, 6, 0, 5, 5, 0, 5, 5, 0, 2, 2, 0, 4, 4, 4,
		4, 0
	);
	-- ��Ŀ 3���滨�����������
	CONSTANT pear : pitch_array3 := (
		-- 1, 1, 1, 1, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 5, 5, 5, 5, 3, 3, 3, 3,
		-- 2, 2, 2, 2, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 0, 3, 3, 3, 3, 5, 5, 5, 5, 3, 3, 3, 3, 2, 2, 2, 2,
		-- 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0

		4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 8, 8, 8, 8, 
		6, 6, 6, 6, 5, 5, 5, 5, 6, 6, 6, 6, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 0, 6, 6, 6, 6, 
		8, 8, 8, 8, 6, 6, 6, 6, 5, 5, 5, 5, 6, 6, 6, 6, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 0, 
		2, 2, 2, 2, 1, 1, 2, 2, 4, 4, 2, 2, 4, 4, 4, 4, 6, 6, 6, 6, 5, 5, 5, 5, 6, 6, 6, 6, 
		5, 5, 5, 5, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 
		4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 8, 8, 8, 8, 6, 6, 6, 6, 5, 5, 5, 5, 6, 6, 6, 6, 
		5, 5, 5, 5, 4, 4, 4, 4, 0, 0, 6, 6, 6, 6, 8, 8, 8, 8, 6, 6, 6, 6, 5, 5, 5, 5, 6, 6, 6, 6,
		5, 5, 5, 5, 4, 4, 4, 4, 0, 0, 2, 2, 2, 2, 1, 1, 2, 2, 4, 4, 2, 2, 4, 4, 4, 4, 6, 6, 6, 6,
		5, 5, 5, 5, 6, 6, 6, 6, 5, 5, 5, 5, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0
	);

	-- 8, 8, 8, 8, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 10, 10, 10, 10, 12, 12, 12, 12, 
	-- 10, 10, 10, 10, 9, 9, 9, 9, 10, 10, 10, 10, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 0, 10, 10, 
	-- 10, 10, 12, 12, 12, 12, 10, 10, 10, 10, 9, 9, 9, 9, 10, 10, 10, 10, 9, 9, 9, 9, 9, 9, 9, 9, 
	-- 8, 8, 8, 8, 0, 0, 6, 6, 6, 6, 5, 5, 6, 6, 8, 8, 6, 6, 8, 8, 8, 8, 10, 10, 10, 10, 
	-- 9, 9, 9, 9, 10, 10, 10, 10, 9, 9 ,9, 9, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 0, 0, 8, 8, 8, 8, 
	-- 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 10, 10, 10, 10, 12, 12, 12, 12, 10, 10, 10, 10, 
	-- 9, 9, 9, 9, 10, 10, 10, 10, 9, 9, 9, 9, 8, 8, 8, 8, 0, 10, 10, 10, 10, 12, 12, 12, 12,
	-- 10, 10, 10, 10, 9, 9, 9, 9, 10, 10, 10, 10, 9, 9, 9, 9, 8, 8, 8, 8, 0 
	-- 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 6, 6, 6, 6, 8, 8, 8, 8, 6, 6, 6, 6,
	-- 5, 5, 5, 5, 6, 6, 6, 6, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 0, 6, 6, 6, 6, 8, 8, 8, 8, 6, 6, 6, 6, 5, 5, 5, 5,
	-- 6, 6, 6, 6, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 0, 0

BEGIN
	-- �����̣����� 8Hz ʱ���źź͵�ǰ��������������
	PROCESS (clk8hz, music_num)
	BEGIN
		-- �����������Ƿ��л�
		IF music_num /= mn_former THEN
			mn_former <= music_num; -- ���¼�¼���������
			ptr1 <= 0; -- �л���Ŀ���ͷ��ʼ����
			ptr2 <= 0;
			ptr3 <= 0;
		ELSE
			-- �� 8Hz ʱ���źŵ������ظ�������ָ��
			IF rising_edge(clk8hz) THEN
				-- ѭ��������Ŀ 1
				IF ptr1 = 239 THEN
					ptr1 <= 0;
				ELSE
					ptr1 <= ptr1 + 1;
				END IF;
				-- ѭ��������Ŀ 2
				IF ptr2 = 181 THEN
					ptr2 <= 0;
				ELSE
					ptr2 <= ptr2 + 1;
				END IF;
				-- ѭ��������Ŀ 3
				IF ptr3 = 255 THEN
					ptr3 <= 0;
				ELSE
					ptr3 <= ptr3 + 1;
				END IF;
			END IF;

			-- ���ݵ�ǰ�������ѡ���������
			CASE music_num IS
				WHEN 0 => -- ��Ŀ 1: С����
					tone2 <= little_star(ptr1);
				WHEN 1 => -- ��Ŀ 2: ��л������
					tone2 <= thx(ptr2);
				WHEN 2 => -- ��Ŀ 3: �滨��
					tone2 <= pear(ptr3);
			END CASE;
		END IF;
	END PROCESS;
END song_arch;